typedef struct packed {
    bit high;
    bit low;
} Dual;
